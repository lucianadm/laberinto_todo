library verilog;
use verilog.vl_types.all;
entity control_motor_vlg_vec_tst is
end control_motor_vlg_vec_tst;
