library verilog;
use verilog.vl_types.all;
entity contador_n_bits_vlg_vec_tst is
end contador_n_bits_vlg_vec_tst;
