library verilog;
use verilog.vl_types.all;
entity decoder4to16_vlg_check_tst is
    port(
        Y0              : in     vl_logic;
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        Y3              : in     vl_logic;
        Y4              : in     vl_logic;
        Y5              : in     vl_logic;
        Y6              : in     vl_logic;
        Y7              : in     vl_logic;
        Y8              : in     vl_logic;
        Y9              : in     vl_logic;
        Y10             : in     vl_logic;
        Y11             : in     vl_logic;
        Y12             : in     vl_logic;
        Y13             : in     vl_logic;
        Y14             : in     vl_logic;
        Y15             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder4to16_vlg_check_tst;
